LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;

ENTITY Processor IS
    PORT (
    );
END ENTITY Processor;

ARCHITECTURE arKAKtectureProcessor OF Processor IS
END ARCHITECTURE arKAKtectureProcessor;